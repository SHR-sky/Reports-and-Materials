module Dram(
    input clk,
    input wb,
    input [4:0] addr,
    input [1:0] lb,
    input [31:0] WriteData,
    input MemWr,

    output reg [31:0] ReadData

);
    //���ݴ洢�����
    reg [31:0] regs[0:31];  //32��32λ�ļĴ���
    always @(addr)begin
       if(wb)begin
            case (lb[1:0])
                2'b00:
                begin
                    if(regs[addr][31] == 1)
                        ReadData <= {24'hffffff, regs[addr][31:24]}; // LB 3:0
                    else if(regs[addr][31] == 0)
                        ReadData <= {24'b0, regs[addr][31:24]}; // LB 3:0
                end
                2'b01: 
                begin
                    if(regs[addr][23] == 1)
                        ReadData <= {24'hffffff, regs[addr][23:16]}; // LB 7:4
                    else if (regs[addr][23] == 0)
                        ReadData <= {24'b0, regs[addr][23:16]}; // LB 7:4
                end
                2'b10: 
                begin
                    if(regs[addr][15] == 1)
                        ReadData <= {24'hffffff, regs[addr][15:8]}; // LB 11:8
                    else if (regs[addr][15] == 0)
                        ReadData <= {24'b0, regs[addr][15:8]}; // LB 11:8
                end
                2'b11: 
                begin
                    if(regs[addr[4:0]][7] == 1)
                        ReadData <= {24'hffffff, regs[addr][7:0]}; // LB 15:12
                    else if (regs[addr[4:0]][7] == 0)
                        ReadData <= {24'b0, regs[addr][7:0]}; // LB 15:12
                end
                default:ReadData <= 0;
            endcase
       end
       else begin
            ReadData = regs[addr];
       end
    end

    //���ݴ洢��д��
    always @(negedge clk) begin
        if(MemWr) regs[addr] = WriteData;
    end

    //���ݴ洢����ʼ��
    integer i;
    initial begin
        for(i=0;i<32;i=i+1) begin
            regs[i] = i*4;
        end
    end
endmodule